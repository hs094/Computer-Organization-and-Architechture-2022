`timescale 1ns / 1 ps
/* ---------------------------------------------------------
*    # COMPUTER ORGANIZATION LABORATORY
*    # AUTUMN SEMESTER 2022
*    # RISC Processor Design
*    # Group No. 60
*    # Abhay Kumar Keshari 20CS10001
*    # Hardik Soni 20CS30023
*---------------------------------------------------------
*/ 
module ALU(
    input signed [31:0] a,
    input signed [31:0] b,
    input ALUsel,
    input [4:0] ALUop,
    output [31:0] result,
    output reg carry,
    output reg sign,
    output reg zero
);

    // Stores carry generated by adder1
    wire carryTemp;
    // Stores 32-bit output of not, adder1, shifter, and, xor, mux1, mux2 respectively from left to right
    wire [31:0]
